-- Libraries required for the operation of the ULA
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


-- Description of the ULA inputs and outputs
entity ULA is

    Port (  clk : in std_logic; -- Clock input 
				button : in std_logic; -- Button input
				switches : in std_logic_vector(3 downto 0); -- Input 4 switches (sw0, sw1, sw2 and sw3)
				leds_out : out std_logic_vector(7 downto 0)); -- Output 8 leds (ld0, ld1, ld2, ld3, ld4, ld5, ld6 and ld7)

end ULA;

-- Description of the ULA behavior
architecture Behavioral of ULA is

	component ULA_debounce -- Incorporate the debounce file
   
	Port(	clk: in std_logic; -- Send clock input
			input: in std_logic; -- Send button input
			debounce: out std_logic); -- Returns debounce pulse
	end component;
	
	component operations is -- Incorporate the operations file
	
	Port(	clk : in std_logic; -- Send clock input
			opcode : in std_logic_vector (2 downto 0); -- Send the operation's code
         A : in std_logic_vector (3 downto 0); -- -- Send the first number inserted
         B : in std_logic_vector (3 downto 0); -- -- Send the second number inserted
			result : out std_logic_vector (7 downto 0)); -- Returns the operation result
	end component;

	-- Signals sent to the operations component
	signal a: std_logic_vector(3 downto 0) := "0000"; -- First number = 0
	signal b: std_logic_vector(3 downto 0) := "0000"; -- Second number = 0
	signal opcode: std_logic_vector(2 downto 0) := "000"; -- Operation = AND
	
	-- Signals returned from the components
	signal result: std_logic_vector(7 downto 0); -- Result of the operation comes from the operations component
	signal debounce: std_logic; -- Debounced pulse comes from the ULA_debounce component

	-- Signals used only in the state machine
	signal leds: std_logic_vector(7 downto 0) := "00000000"; -- Displays output = 0
	signal state: std_logic_vector(1 downto 0) := "00"; -- Controls the state of the state machine, initial state 0
	
begin

-- DUT of debounce, links the signals of this file with the inputs and outputs of the debounce component
	deb_dut: ULA_debounce port map (
        clk      => clk,
        input    => button,
        debounce => debounce
    );

-- DUT of operations, links the signals of this file with the inputs and outputs of the operations component	 
	 op_dut: operations port map (
        clk    => clk,
		  opcode => opcode,
        a      => A,
        b      => B,
		  result => result
    );
	 
-- Links the signal with what should be displayed on the LEDs using the LED pins (outputs should be assigned outside the process)
	leds_out <= leds;
 
-- Clock-dependent sequential process with the state machine
process(clk)

	--It needs to have an operation variable to make the decision to jump states within the same clock cycle
	variable operation_var : std_logic_vector(2 downto 0); -- Chosen operation variable
	
begin
	if (clk'event and clk = '1') then -- On the rising edge of the clock
    	if (debounce = '1') then -- On the debounced pulse
			
			case state is -- According to the current state
			
				when "00" => -- When state is 00, register the chosen operation
				
					-- Links the switch inputs with what should be displayed on the LEDs and with the operation variable
					for i in 0 to 2 loop
						operation_var(i) := switches(i);
						leds(i) <= switches(i);
					end loop;
					
					-- Pads the most significant LEDs with zero
					for i in 0 to 4 loop
						leds(3+i) <= '0';
					end loop;
					
					-- If the operation is modulo, skip one state
					if (operation_var = "011") then
						state <= "11";
					else
						state <= "01";
					end if;
					
					-- The chosen operation signal is linked to the operation variable
					opcode <= operation_var;

				
				when "01" => -- When the state is 01, register the first number
				
					a <= "0000"; -- Ensures that the number is zeroed
				
					-- Links the switch inputs with what should be displayed on the LEDs and with the first number signal
					for i in 0 to 3 loop
						a(i) <= switches(i);
						leds(i) <= switches(i);
					end loop;
					
					-- Pads the most significant LEDs with zero
					for i in 0 to 3 loop
						leds(4+i) <= '0';
					end loop;
					
					-- Changes to the next state
					state <= "11";

					
				when "11" => -- When the state is 11, register the second number
				
					b <= "0000"; -- Ensures that the number is zeroed
				
					-- Links the switch inputs with what should be displayed on the LEDs and with the second number signal
					for i in 0 to 3 loop
						b(i) <= switches(i);
						leds(i) <= switches(i);
					end loop;
					
					-- Pads the most significant LEDs with zero
					for i in 0 to 3 loop
						leds(4+i) <= '0';
					end loop;
					
					-- Changes to the next state
					state <= "10";
				
				when "10" => -- When the state is 10, it should display/register the result
					
					leds <= result; -- The result returned from the operations file should be displayed on the LEDs
					state <= "00"; -- Changes to the first state
				
				when others => -- In case of error
					leds <= "00000000";
					state <= "00";
					
			end case;
		end if;
	end if;
end process;

end Behavioral; 
